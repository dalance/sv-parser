`define A \
  initial begin // comment \
  end

module test();

initial begin
  end

endmodule
