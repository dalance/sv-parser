// First comment
`default_nettype none
// Middle comment
`resetall
// Last comment
