class test21 extends base_class /* base class*/;
	int a;
	int b;
	function int funcname();
		return 2;
	endfunction : funcname
endclass : test21