
`define A(a)
`A // Macro called without required argument.

