`define MOD_INST u_mysubmod
module mymod;
mysubmod `MOD_INST ();
endmodule
