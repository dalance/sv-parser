// In the next comment, there are non-UTF8 bytes.
module M;
// Non-UTF8:X������X
endmodule
