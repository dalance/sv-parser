
`A // Macro called without definition.

