`define A \
  initial begin // comment \
  end

module test();

`A

endmodule
