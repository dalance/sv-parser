module a;
initial begin
    if (3 == 0) begin
    end
end
endmodule
