/*
The compiler directives described in this annex are for informative purposes only and are not part of this
standard.
This annex describes additional compiler directives as companions to the compiler directives described in
Clause 22. The compiler directives described in this annex may not be available in all implementations of
SystemVerilog. The following compiler directives are described in this annex:
*/


`delay_mode_distributed //[E.4]
`delay_mode_path //[E.5]
