module and_op (a, b, c);
`include "test2.svh" endmodule
