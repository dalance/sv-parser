module a;
reg \`~!-_=+\|[]{};:'"",./<>?  ;
endmodule
