`define NAME 42 // Comment
interface foo #(WIDTH = `NAME) ();
endinterface
