module a;
initial begin
    if (`__LINE__ == 0) begin
    end
end
endmodule
