module and_op (a, b, c);
output a;
input b, c;

wire a = b & c;

endmodule
