module and_op (a, b, c);
  // a
  `include "test2.svh"
endmodule
