module and_op (a, b, c);
`include "test3.sv"
endmodule
