`define A 42 // Comment
interface i #(p = 42) (); endinterface
