module and_op (a, b, c);
output a;
input b, c;

and a1 (a,b,c);

endmodule
