//top
`resetall
`timescale 10 us / 100 ns
`default_nettype wire
//first
`default_nettype none//middle
//last
`unconnected_drive pull0
`unconnected_drive pull1
`nounconnected_drive
`celldefine
`endcelldefine
`pragma foo
`pragma foo bar
`line 5 "foo" 0
`begin_keywords "1800-2017"
`end_keywords
