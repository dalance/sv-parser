`define A 42 // Comment
interface i #(p = `A) (); endinterface
