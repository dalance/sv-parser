`define a `a
// direct recursion
`a
