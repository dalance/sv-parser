module a;
`define A "aaa"
`define \B "bbb"
initial begin
$display("aaa");
$display("aaa");
$display("bbb");
$display("bbb");
end
endmodule
