// __FILE__ = `__FILE__

// This block SHOULD be emitted from the preprocessor.


// Emitted instead.


// The following define should have no effect.
`define __FILE__ "FOO"

// The following undef should have no effect.
`undef __FILE__

// NOTE: Comparison against expected value are destined to fail in testcase.
