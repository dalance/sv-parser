`define MOD_INST u_mysubmod
module mymod;
mysubmod u_mysubmod() ;
endmodule
